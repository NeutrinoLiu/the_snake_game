module vga(clk,
	//map,
			snake_x,
			snake_y,
			apple_x,
			apple_y,

	RGB,hs,vs,blank,sync,clk25);
input clk;
//input [64*48-1:0] map;

input [599:0] snake_x, snake_y;
input [29:0] apple_x, apple_y;




output[24:1] RGB;
output clk25;
output sync;
reg sync=0;
reg[24:1] RGB=000000;
output vs,hs,blank;
reg vs,hs,blank;
reg [5:0] x=0, y=0;

reg[9:0] cntv=0;
reg[9:0] cnth=0;
reg clk25=1'b0;

always@(posedge clk)
	begin
		clk25=~clk25;
	end

always@(posedge clk25)
	begin
		if(cnth==799)
			begin
				cnth=0;
				if(cntv==524)cntv=0;
				else cntv=cntv+1;
			end
		else cnth=cnth+1;
	end

always@(posedge clk)
	begin
		if(cnth<96)hs=1'b0;
		else hs=1'b1;

		if(cntv<2)vs=1'b0;
		else vs=1'b1;
	end	

always @(posedge clk)
	begin
		if(cntv<35||cntv>514||cnth<144||cnth>783) blank=1'b0;
		else blank=1'b1;
	end

wire answer;
inquiry q1(
			snake_x,
			snake_y,
			apple_x,
			apple_y,
			x,
			y,
			answer
			);

always @( x or y or answer)
	begin
		if (answer) RGB = 24'hffffff;
		else RGB = 24'h000000;
	end

always @(cntv or cnth)
begin
	case (cntv)
35,36,37,38,39,40,41,42,43,44: y = 0;
45,46,47,48,49,50,51,52,53,54: y = 1;
55,56,57,58,59,60,61,62,63,64: y = 2;
65,66,67,68,69,70,71,72,73,74: y = 3;
75,76,77,78,79,80,81,82,83,84: y = 4;
85,86,87,88,89,90,91,92,93,94: y = 5;
95,96,97,98,99,100,101,102,103,104: y = 6;
105,106,107,108,109,110,111,112,113,114: y = 7;
115,116,117,118,119,120,121,122,123,124: y = 8;
125,126,127,128,129,130,131,132,133,134: y = 9;
135,136,137,138,139,140,141,142,143,144: y = 10;
145,146,147,148,149,150,151,152,153,154: y = 11;
155,156,157,158,159,160,161,162,163,164: y = 12;
165,166,167,168,169,170,171,172,173,174: y = 13;
175,176,177,178,179,180,181,182,183,184: y = 14;
185,186,187,188,189,190,191,192,193,194: y = 15;
195,196,197,198,199,200,201,202,203,204: y = 16;
205,206,207,208,209,210,211,212,213,214: y = 17;
215,216,217,218,219,220,221,222,223,224: y = 18;
225,226,227,228,229,230,231,232,233,234: y = 19;
235,236,237,238,239,240,241,242,243,244: y = 20;
245,246,247,248,249,250,251,252,253,254: y = 21;
255,256,257,258,259,260,261,262,263,264: y = 22;
265,266,267,268,269,270,271,272,273,274: y = 23;
275,276,277,278,279,280,281,282,283,284: y = 24;
285,286,287,288,289,290,291,292,293,294: y = 25;
295,296,297,298,299,300,301,302,303,304: y = 26;
305,306,307,308,309,310,311,312,313,314: y = 27;
315,316,317,318,319,320,321,322,323,324: y = 28;
325,326,327,328,329,330,331,332,333,334: y = 29;
335,336,337,338,339,340,341,342,343,344: y = 30;
345,346,347,348,349,350,351,352,353,354: y = 31;
355,356,357,358,359,360,361,362,363,364: y = 32;
365,366,367,368,369,370,371,372,373,374: y = 33;
375,376,377,378,379,380,381,382,383,384: y = 34;
385,386,387,388,389,390,391,392,393,394: y = 35;
395,396,397,398,399,400,401,402,403,404: y = 36;
405,406,407,408,409,410,411,412,413,414: y = 37;
415,416,417,418,419,420,421,422,423,424: y = 38;
425,426,427,428,429,430,431,432,433,434: y = 39;
435,436,437,438,439,440,441,442,443,444: y = 40;
445,446,447,448,449,450,451,452,453,454: y = 41;
455,456,457,458,459,460,461,462,463,464: y = 42;
465,466,467,468,469,470,471,472,473,474: y = 43;
475,476,477,478,479,480,481,482,483,484: y = 44;
485,486,487,488,489,490,491,492,493,494: y = 45;
495,496,497,498,499,500,501,502,503,504: y = 46;
505,506,507,508,509,510,511,512,513,514: y = 47;
default: y = 0;
endcase

	case (cnth)
144,145,146,147,148,149,150,151,152,153: x = 0;
154,155,156,157,158,159,160,161,162,163: x = 1;
164,165,166,167,168,169,170,171,172,173: x = 2;
174,175,176,177,178,179,180,181,182,183: x = 3;
184,185,186,187,188,189,190,191,192,193: x = 4;
194,195,196,197,198,199,200,201,202,203: x = 5;
204,205,206,207,208,209,210,211,212,213: x = 6;
214,215,216,217,218,219,220,221,222,223: x = 7;
224,225,226,227,228,229,230,231,232,233: x = 8;
234,235,236,237,238,239,240,241,242,243: x = 9;
244,245,246,247,248,249,250,251,252,253: x = 10;
254,255,256,257,258,259,260,261,262,263: x = 11;
264,265,266,267,268,269,270,271,272,273: x = 12;
274,275,276,277,278,279,280,281,282,283: x = 13;
284,285,286,287,288,289,290,291,292,293: x = 14;
294,295,296,297,298,299,300,301,302,303: x = 15;
304,305,306,307,308,309,310,311,312,313: x = 16;
314,315,316,317,318,319,320,321,322,323: x = 17;
324,325,326,327,328,329,330,331,332,333: x = 18;
334,335,336,337,338,339,340,341,342,343: x = 19;
344,345,346,347,348,349,350,351,352,353: x = 20;
354,355,356,357,358,359,360,361,362,363: x = 21;
364,365,366,367,368,369,370,371,372,373: x = 22;
374,375,376,377,378,379,380,381,382,383: x = 23;
384,385,386,387,388,389,390,391,392,393: x = 24;
394,395,396,397,398,399,400,401,402,403: x = 25;
404,405,406,407,408,409,410,411,412,413: x = 26;
414,415,416,417,418,419,420,421,422,423: x = 27;
424,425,426,427,428,429,430,431,432,433: x = 28;
434,435,436,437,438,439,440,441,442,443: x = 29;
444,445,446,447,448,449,450,451,452,453: x = 30;
454,455,456,457,458,459,460,461,462,463: x = 31;
464,465,466,467,468,469,470,471,472,473: x = 32;
474,475,476,477,478,479,480,481,482,483: x = 33;
484,485,486,487,488,489,490,491,492,493: x = 34;
494,495,496,497,498,499,500,501,502,503: x = 35;
504,505,506,507,508,509,510,511,512,513: x = 36;
514,515,516,517,518,519,520,521,522,523: x = 37;
524,525,526,527,528,529,530,531,532,533: x = 38;
534,535,536,537,538,539,540,541,542,543: x = 39;
544,545,546,547,548,549,550,551,552,553: x = 40;
554,555,556,557,558,559,560,561,562,563: x = 41;
564,565,566,567,568,569,570,571,572,573: x = 42;
574,575,576,577,578,579,580,581,582,583: x = 43;
584,585,586,587,588,589,590,591,592,593: x = 44;
594,595,596,597,598,599,600,601,602,603: x = 45;
604,605,606,607,608,609,610,611,612,613: x = 46;
614,615,616,617,618,619,620,621,622,623: x = 47;
624,625,626,627,628,629,630,631,632,633: x = 48;
634,635,636,637,638,639,640,641,642,643: x = 49;
644,645,646,647,648,649,650,651,652,653: x = 50;
654,655,656,657,658,659,660,661,662,663: x = 51;
664,665,666,667,668,669,670,671,672,673: x = 52;
674,675,676,677,678,679,680,681,682,683: x = 53;
684,685,686,687,688,689,690,691,692,693: x = 54;
694,695,696,697,698,699,700,701,702,703: x = 55;
704,705,706,707,708,709,710,711,712,713: x = 56;
714,715,716,717,718,719,720,721,722,723: x = 57;
724,725,726,727,728,729,730,731,732,733: x = 58;
734,735,736,737,738,739,740,741,742,743: x = 59;
744,745,746,747,748,749,750,751,752,753: x = 60;
754,755,756,757,758,759,760,761,762,763: x = 61;
764,765,766,767,768,769,770,771,772,773: x = 62;
774,775,776,777,778,779,780,781,782,783: x = 63;
default: x = 0;
endcase

end


endmodule
